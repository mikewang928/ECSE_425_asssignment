library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fetch is

port(
	instruction : out std_logic_vector(31 downto 0);
);
end fetch;

architecture arch of fetch is


begin



end arch;