library ieee;

use ieee.std_logic_1164.all; -- allows use of the std_logic_vector type
use ieee.numeric_std.all; -- allows use of the unsigned type

PACKAGE memory_constants IS

	constant dm_depth : integer := 65536;

END memory_constants;
