library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity execution is
	port(
		clk : in std_logic;
		
	);
end execution;

architecture arch of execution is



begin



end arch;